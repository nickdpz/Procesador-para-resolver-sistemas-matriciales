use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use IEEE.numeric_std.all;

entity Prueba is
end Prueba;

architecture Behavioral of Prueba is

begin


end Behavioral;

